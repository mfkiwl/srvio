/*
* <decode.svh>
* 
* Copyright (c) 2021 Yosuke Ide <yosuke.ide@keio.jp>
* 
* This software is released under the MIT License.
* https://opensource.org/licenses/mit-license.php
*/

`ifndef _DECODE_SVH_INCLUDED_
`define _DECODE_SVH_INCLUDED_

//***** Functional Unit configuration
typedef struct {
};


typedef struct {
} Decode_t;

`endif //_DECODE_SVH_INCLUDED_
