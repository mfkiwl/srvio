/*
* <io_config.vh>
*
* Copyright (c) 2021 Yosuke Ide <yosuke.ide@keio.jp>
*
* This software is released under the MIT License.
* https://opensource.org/licenses/mit-license.php
*/

`ifndef _IO_CONFIG_H_INCLUDED_
`define _IO_CONFIG_H_INCLUDED_

// 吾輩はio_config.hである。中身はまだない。

`endif
