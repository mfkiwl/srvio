/*
* <complex_dec.sv>
* 
* Copyright (c) 2021 Yosuke Ide <yosuke.ide@keio.jp>
* 
* This software is released under the MIT License.
* https://opensource.org/licenses/mit-license.php
*/

`include "stddef.vh"
`include "cpu_config.svh"

module complex_dec #(
	parameter ADDR = `AddrWidth,
	parameter DATA = `DataWidth
)(
);

endmodule
