/*
* <config.vh>
*
* Copyright (c) 2021 Yosuke Ide <yosuke.ide@keio.jp>
*
* This software is released under the MIT License.
* https://opensource.org/licenses/mit-license.php
*/

`ifndef _CONFIG_SVH_INCLUED_
`define _CONFIG_SVH_INCLUDED_

`include "process_config.svh"
`include "cpu_config.svh"
`include "io_config.svh"

//**** TODO: concat all configs

`endif //_CONFIG_SVH_INCLUED_
